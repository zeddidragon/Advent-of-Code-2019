module main

import advent

fn main() {
  advent.code()
}
