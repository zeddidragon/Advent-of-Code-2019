module advent

pub fn code() {
  day01()
}
