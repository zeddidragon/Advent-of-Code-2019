module advent

fn day(d int, part int) {
  println("Day $d - $part")
  println("===========")
}

fn max(a int, b int) int {
  if(a > b) { return a }
  return b
}

fn arr_copy(arr []int) []int {
  return arr.map(it)
}
