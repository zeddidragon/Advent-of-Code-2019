module advent

pub fn code() {
  day01()
  day02()
  day03()
  day04()
}
