module advent

pub fn code() {
  day01()
  day02()
}
