module advent

pub fn day18() {
	println('I give up')
}
